module adv7393_debug #(parameter DEBUG_ENA = 0) (
  input  clk    ,
  input  rst    ,
  input  clk_pix,
  output invalid
);





endmodule
